//
// Register
//
// Hardik Sharma
// (hsharma@gatech.edu)

/*
module sum:
  wire(int)-reg-wire(out)
  a register with sync;
功能,用于做delay时序赋值(只能delay半个周期,即一个下降沿或者上升沿),或者存储数据
*/

`timescale 1ns/1ps
module register_sync #(
  parameter integer WIDTH                 = 8
) (
  input  wire                             clk,
  input  wire                             reset,
  // input  wire                             enable,
  input  wire        [ WIDTH -1 : 0 ]     in,
  output wire        [ WIDTH -1 : 0 ]     out
);

  reg [ WIDTH -1 : 0 ] out_reg;//internal reg 

  always @(posedge clk)//sync clock
  begin
    // if (reset)
      // out_reg <= 'b0;
    // else if (enable)
      out_reg <= in;
  end

  assign out = out_reg;

endmodule
